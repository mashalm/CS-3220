module EggTimerController();