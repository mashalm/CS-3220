library verilog;
use verilog.vl_types.all;
entity TimerController_testbench is
end TimerController_testbench;
